library verilog;
use verilog.vl_types.all;
entity tf_button is
end tf_button;
