library verilog;
use verilog.vl_types.all;
entity tf_relays is
end tf_relays;
