library verilog;
use verilog.vl_types.all;
entity tf_adc is
end tf_adc;
